interface intf(input logic clk);
    logic d, q, q_inverted;
endinterface:intf